Testddddsdsddsdad
eweaweawe
Editesewsrdsadssadsadssdasdsadsadd
ssdasddsdsadsdfdsf
dsdssadasdasdsad
My mind!! Twestese wewessdsaddsaddsadasdsadasdasddsadas sadasd
Omg this is so cool


Other way test