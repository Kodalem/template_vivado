-- THIS IS A DUMMY FILE FOR DESIGN SOURCES