-- THIS IS A DUMMYsdsasdsa FILaaaaaaE FORdasds SIMULATION SOURCES