-- THIS IS A DUMMY FILE FOR SIMULATION SOURCES